`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 31.10.2021 00:39:28
// Design Name: 
// Module Name: alufirst
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module alufirst(
   input [5:0] x1,y1,
   output [5:0] c1
    );
   assign c1 = x1;  //we want the output A
endmodule
