module alusecond(
   input [5:0] x2,y2,
   output [5:0] c2
    );
   assign c2 = y2; //we want the output B
endmodule